.title KiCad schematic
C1 + NC_01 CP1
R1 + + R_US
.end
